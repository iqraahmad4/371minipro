module main(col,row/*,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7*/);
input[3:0] col;
input[3:0]row;
//GetRowAndCol(); //see which button has been pressed
//CheckTypeAndStore(row, col); //function that checks what button has been pressed if its an integer or an operation
					//if number make sure doesnt exceed 8 digits(maybe) and store digit store. No more than 8 digits can be stored at a time
					//allow indicator to see i a number is negatie need special case for detecting negative. 
					//Dont count negative as an operation if at beginning iof a number and after a previous opration has ben pressed
					//if operation store which operation has been pressed
					//store all digits after operator has been pressed in a second container
//if(row== && col==)
					//begin calculation after equal hass been pressed
					//to begin operation  go to the corresponding function to the operatiion
					//take the two numbers stored if bigger than 8 digits display nothing
					//add to numbers create case for negatives 
					//display numbers then clear
//DisplayAns();					//display sum
					
endmodule